module and_4bit(out,in1,in2);
input [3:0] in1, in2;
output [3:0] out;

and t1(out[3], in1[3], in2[3]);
and t2(out[2], in1[2], in2[2]);
and t3(out[1], in1[1], in2[1]);
and t4(out[0], in1[0], in2[0]);
	 
endmodule